module FullAdder(a,b,c,o1,o2);
input a,b,c;
output o1,o2;
wire d,e,f;
xor x1(d,b,c);
xor x2(o1,d,a);
and A1(e,d,a);
and A2(f,b,c);
or or1(o2,e,f);
endmodule


module four_bit_adder(a,b,o);
input[3:0] a;
input[3:0] b;
output[3:0] o;
reg t;
always t=0;
reg[3:0] c;
FullAdder F1(a[0],b[0],t,o[0],c[0]);
FullAdder F2(a[1],b[1],c[0],o[1],c[1]);
FullAdder F3(a[2],b[2],c[1],o[2],c[2]);
Fulladder F4(a[3],b[3],c[2],o[3],c[3]);
endmodule


module four_bit_sub(a,b,o);
input[3:0] a;
input[3:0] b;
output[4:0] o;
reg[3:0] c;
always@(b) c=b^1;
wire[4:0] d;
reg[3:0] e;
always e[0]=1;
always e[1]=0;
always e[2]=0;
always e[3]=0;
four_bit_adder f1(c,e,d);
four_bit_adder f2(a,d,o);
endmodule


module four_bit_comp(a0,a1,a2,a3,b0,b1,b2,b3,o1,o2,o3);
input a0,a1,a2,a3;
input b0,b1,b2,b3;
inout o1,o2,o3;
wire s1,s2,s3,s4,s5,s6,s7,s8,p,q,b01,b11,b21,b31,o;
not N0(b01,b0);
not N1(b11,b1);
not N2(b21,b2);
not N3(b31,b3);
and A1(s1,a3,b3);
and A2(s2,a2,b21,s5);
and A3(s3,a1,b11,s5,s6);
and A4(s4,a0,b01,s5,s6,s7);
or R1(p,s1,s2,s3,s4);
not N4(o,p);
xor X3(s5,a3,b3);
xor X2(s6,a2,b2);
xor X1(s7,a1,b1);
xor X0(s8,a0,b0);
and(q,s5,s6,s7,s8);
not N5(o3,q);
or R2(o2,o3,o1);
endmodule


module gcd_cal (A,B,C);
input [3:0] A,B;
output [3:0] C;
wire [4:0]sub;

reg [7:0] p;
wire AgB,BgA,AeB;
wire m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,m15,m16;
wire ns0,ns1,ns2,ns3,check,nBgA;
four_bit_comp f1(A[0],A[1],A[2],A[3],B[0],B[1],B[2],B[3],AgB,BgA,AeB);
not n0(nBgA,BgA);
and s1(m1,A[0],nBgA);
and s2(m2,A[0],BgA);
and s3(m3,A[1],nBgA);
and s4(m4,A[1],BgA);
and s5(m5,A[2],nBgA);
and s6(m6,A[2],BgA);
and s7(m7,A[3],nBgA);
and s8(m8,A[3],BgA);
and s9(m9,B[0],nBgA);
and s10(m10,B[0],BgA);
and s11(m11,B[1],nBgA);
and s12(m12,B[1],BgA);
and s13(m13,B[2],nBgA);
and s14(m14,B[2],BgA);
and s15(m15,B[3],nBgA);
and s16(m16,B[3],BgA);
or  q1(p[0],m1,m2);
or  q2(p[1],m3,m4);
or  q3(p[2],m5,m6);
or  q4(p[3],m7,m8);
or  q5(p[4],m9,m10);
or  q6(p[5],m11,m12);
or  q7(p[6],m13,m14);
or  q8(p[7],m15,m16);
assign A[3:0]=p[3:0];
assign B[3:0]=p[7:4];

four_bit_sub f2(A[3:0],B[3:0],sub[4:0]);
not n1(ns0,sub[0]);
not n2(ns1,sub[1]);
not n3(ns2,sub[2]);
not n4(ns3,sub[3]);
and w1(C[0],ns0,B[0]);
and w2(C[1],ns1,B[1]);
and w3(C[2],ns2,B[2]);
and w4(C[3],ns3,B[3]);

nand a1(check,ns0,ns1,ns2,ns3);//check is 0 when sub is 0000,else check is 1
and a2(A[0],check,sub[0]);
and a3(A[1],check,sub[1]);
and a4(A[2],check,sub[2]);
and a5(A[3],check,sub[3]);

and a6(B[0],check,p[4]);
and a7(B[1],check,p[5]);
and a8(B[2],check,p[6]);
and a9(B[3],check,p[7]);

endmodule
